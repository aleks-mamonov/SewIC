.subckt p_mos S D
* Subcircuit Body
.ends p_mos